// 4 bit ripple carry adder
// http://fullchipdesign.com/fulladder.htm
// http://fullchipdesign.com/4_bit_binary_adder.htm

module half_adder(S,C,x,y);
    output S,C;
    input x,y;
    
endmodule
