// 8 to 1 multiplexer
// https://www.electronicshub.org/multiplexerandmultiplexing/#8-to-1_Multiplexer

module multiplexer_8_to_1(Y,D,S);
    output Y;
    input [0:7] D;
    input [0:2] S;
    wire [0:2] not_S;
    wire [0:7] I;
    not G1(not_S[0],S[0]);
    not G2(not_S[1],S[1]);
    not G3(not_S[2],S[2]);
    and G4(I[0],D[0],not_S[0],not_S[1],not_S[2]);
    and G5(I[1],D[1],S[0],not_S[1],not_S[2]);
    and G6(I[2],D[2],not_S[0],S[1],not_S[2]);
    and G7(I[3],D[3],S[0],S[1],not_S[2]);
    and G8(I[4],D[4],not_S[0],not_S[1],S[2]);
    and G9(I[5],D[5],S[0],not_S[1],S[2]);
    and G10(I[6],D[6],not_S[0],S[1],S[2]);
    and G11(I[7],D[7],S[0],S[1],S[2]);
    or G12(Y,I[0],I[2],I[3],I[4],I[5],I[6],I[7]);
endmodule

module test_multiplexer_8_to_1();
    wire Y;
    reg [0:7] D;
    reg [0:2] S;
    multiplexer_8_to_1 G(Y,D,S);
    initial 
	begin
	    D=8'b10101011;
	    #50 S=4'b000;
	    #50 S=4'b100;
	    #50 S=4'b010;
	    #50 S=4'b110;
	    #50 S=4'b001;
	    #50 S=4'b101;
	    #50 S=4'b011;
	    #50 S=4'b111;
	end
endmodule
